LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY REG_DCC_TB IS
END ENTITY;

ARCHITECTURE tb OF REG_DCC_TB IS
  COMPONENT REG_DCC
    PORT (
      clk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      load : IN STD_LOGIC;
      shift : IN STD_LOGIC;
      read : IN STD_LOGIC;
      trame_in : IN STD_LOGIC_VECTOR(41 DOWNTO 0);
      emptyy : OUT STD_LOGIC;
      decale : OUT STD_LOGIC;
      data_bit : OUT STD_LOGIC
    );
  END COMPONENT;

  SIGNAL clk : STD_LOGIC;
  SIGNAL reset : STD_LOGIC;
  SIGNAL load : STD_LOGIC;
  SIGNAL shift : STD_LOGIC;
  SIGNAL read : STD_LOGIC;
  SIGNAL trame_in : STD_LOGIC_VECTOR(41 DOWNTO 0);
  SIGNAL emptyy : STD_LOGIC;
  SIGNAL decale : STD_LOGIC;
  SIGNAL data_bit : STD_LOGIC;
  --constant clk_period : time := 1000ns; 

  TYPE tbsigs IS RECORD
    clk : STD_LOGIC;
    reset : STD_LOGIC;
    load : STD_LOGIC;
    shift : STD_LOGIC;
    read : STD_LOGIC;
    trame_in : STD_LOGIC_VECTOR(41 DOWNTO 0);
  END RECORD;

  TYPE testv IS ARRAY (NATURAL RANGE <>) OF tbsigs;
  CONSTANT tv : testv :=(
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '1', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '1', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '1', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '1', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '1', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '1', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '1', '1', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '1', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010"),
  ('0', '0', '0', '0', '0', "101010101010101010101010101010101010101010"), ('1', '0', '0', '0', '0', "101010101010101010101010101010101010101010")
  );

BEGIN
instance : REG_DCC PORT MAP(clk => clk, reset => reset, load => load, shift => shift, read => read, trame_in => trame_in, emptyy => emptyy, decale => decale, data_bit => data_bit);
clocking : PROCESS
VARIABLE vtv : tbsigs;
  BEGIN
    FOR i IN tv'RANGE LOOP
      vtv := tv(i);
      reset <= vtv.reset;
      clk <= vtv.clk;
      load <= vtv.load;
      shift <= vtv.shift;
      read <= vtv.read;
      trame_in <= vtv.trame_in;
      WAIT FOR 5 ns;
    END LOOP;
    WAIT;
  END PROCESS clocking;
END TB;