LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY MAE_TB IS
END ENTITY;
ARCHITECTURE tb OF MAE_TB IS

  COMPONENT mae

    PORT (
      clk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      
      --from REG
      emptyFreg : IN STD_LOGIC;
      bitFreg : IN STD_LOGIC;
      shiftedFreg : IN STD_LOGIC;
      
      --from zero
      startedFzero : IN STD_LOGIC;
      endFzero : IN STD_LOGIC;

      --from zero
      startedFone : IN STD_LOGIC;
      endFone : IN STD_LOGIC;

      --from tempo
      endFtempo : IN STD_LOGIC;

      --OUTPUTS  
      --reset the system
      rst_sys : OUT STD_LOGIC;

      -- to reg
      load2reg : OUT STD_LOGIC;
      shift2reg : OUT STD_LOGIC;
      read2reg : OUT STD_LOGIC;

      --to send_zero_one modules
      enable2one : OUT STD_LOGIC;
      enable2zero : OUT STD_LOGIC;
      
      --to tempo
      enable2tempo : OUT STD_LOGIC
    );
  END COMPONENT;

  SIGNAL clk : STD_LOGIC;
  SIGNAL reset : STD_LOGIC;
  SIGNAL emptyFreg : STD_LOGIC;
  SIGNAL bitFreg : STD_LOGIC;
  SIGNAL shiftedFreg : STD_LOGIC;
  SIGNAL startedFzero : STD_LOGIC;
  SIGNAL endFzero : STD_LOGIC;
  SIGNAL startedFone : STD_LOGIC;
  SIGNAL endFone : STD_LOGIC;
  SIGNAL endFtempo : STD_LOGIC;
  SIGNAL rst_sys : STD_LOGIC;
  SIGNAL load2reg : STD_LOGIC;
  SIGNAL shift2reg : STD_LOGIC;
  SIGNAL read2reg : STD_LOGIC;
  SIGNAL enable2one : STD_LOGIC;
  SIGNAL enable2zero : STD_LOGIC;

  SIGNAL enable2tempo : STD_LOGIC;
  --constant clk_period : time := 1000ns; 
  TYPE tbsigs IS RECORD
    clk : STD_LOGIC;
    reset : STD_LOGIC;
    emptyFreg : STD_LOGIC;
    bitFreg : STD_LOGIC;
    shiftedFreg : STD_LOGIC;
    startedFzero : STD_LOGIC;
    endFzero : STD_LOGIC;
    startedFone : STD_LOGIC;
    endFone : STD_LOGIC;
    endFtempo : STD_LOGIC;
  END RECORD;

  TYPE testv IS ARRAY (NATURAL RANGE <>) OF tbsigs;
  CONSTANT tv : testv :=
  (
  ('0', '1', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), --1
  ('0', '1', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), --2
  ('0', '1', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --3
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '1'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '1'), --4
  ('0', '0', '1', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '1', '0', '0', '0', '0', '0', '0', '0'), --5
  ('0', '0', '1', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '1', '0', '0', '0', '0', '0', '0', '0'), --6
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --7
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --8
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --9
  ('0', '0', '0', '0', '0', '1', '1', '0', '0', '0'), ('1', '0', '0', '0', '0', '1', '1', '0', '0', '0'), --10
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --11
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --12
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --13
  ('0', '0', '0', '0', '1', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '1', '0', '0', '0', '0', '0'), --14
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --15
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --16
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --17
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --18
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --19
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --20
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --21
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --22    
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --23
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --24
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --25
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --26
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --27
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --28
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --29
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --30
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --31
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --32
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --33
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --34
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --35
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --36
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --37
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --38
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --39
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --40
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --41
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --42
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), --43
  ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), ('1', '0', '0', '0', '0', '0', '0', '0', '0', '0') --44  
  );

BEGIN
INSTANCE : mae
  PORT MAP(
    clk => clk, reset => reset, emptyFreg => emptyFreg, bitFreg => bitFreg, shiftedFreg => shiftedFreg, startedFzero => startedFzero, endFzero => endFzero, startedFone => startedFone, endFone => endFone, endFtempo => endFtempo, rst_sys => rst_sys, load2reg => load2reg, shift2reg => shift2reg,
    read2reg => read2reg, enable2one => enable2one, enable2zero => enable2zero, enable2tempo => enable2tempo);

clocking : PROCESS
  VARIABLE vtv : tbsigs;
  BEGIN
    FOR i IN tv'RANGE LOOP
      vtv := tv(i);
      reset <= vtv.reset;
      clk <= vtv.clk;
      emptyFreg <= vtv.emptyFreg;
      bitFreg <= vtv.bitFreg;
      shiftedFreg <= vtv.shiftedFreg;
      startedFzero <= vtv.startedFzero;
      endFzero <= vtv.endFzero;
      startedFone <= vtv.startedFone;
      endFone <= vtv.endFone;
      endFtempo <= vtv.endFtempo;
      WAIT FOR 5 ns;
    END LOOP;
    WAIT;
END PROCESS clocking;
END TB;